library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity mux_16x1_8bit is
    port (
        inputs   : in  STD_LOGIC_VECTOR(127 downto 0); -- 16 inputs, each 8-bit wide
        sel      : in  STD_LOGIC_VECTOR(15 downto 0); -- 16-bit 1-hot select signal
        sel_4bit : in  std_logic_vector(3 downto 0);
        output   : out STD_LOGIC_VECTOR(7 downto 0) -- 8-bit output
    );
end entity mux_16x1_8bit;

architecture Structural of mux_16x1_8bit is

    -- Declare the 2x1 8-bit multiplexer component
    component mux_16x1 is
        port (
            inputs      : in  STD_LOGIC_VECTOR(15 downto 0); -- 16-bit input vector
            sel         : in  STD_LOGIC_VECTOR(3 downto 0);  -- 4-bit select signal
            sel_one_hot : in  std_logic_vector(15 downto 0);
            output      : out STD_LOGIC                      -- Output of the multiplexer
        );
    end component mux_16x1;

    signal bits : std_logic_vector(127 downto 0);

begin

    gen_1: for i in 0 to 7 generate
        bits((16 * (i + 1) - 1) downto (16 * i)) <=
            (
                inputs(i + 120),
                inputs(i + 112),
                inputs(i + 104),
                inputs(i + 96),
                inputs(i + 88),
                inputs(i + 80),
                inputs(i + 72),
                inputs(i + 64),
                inputs(i + 56),
                inputs(i + 48),
                inputs(i + 40),
                inputs(i + 32),
                inputs(i + 24),
                inputs(i + 16),
                inputs(i + 8),
                inputs(i)
            );
    end generate;

    gen_2: for i in 0 to 7 generate
        select_out: entity work.mux_16x1(Structural)
        port map (
            inputs      => bits(127 - (16 * i) downto 127 - (16 * i) - 15),
            sel         => sel_4bit,
            sel_one_hot => sel,
            output      => output(7 - i)
        );
    end generate;

end architecture Structural;
