-- Created by @(#)$CDS: vhdlin version 6.1.8-64b 06/22/2022 16:17 (sjfhw317) $
-- on Tue Dec  3 11:52:04 2024


architecture Structural of or_2x1 is

begin
    output <= A or B;

end Structural;
