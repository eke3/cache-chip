-- Created by @(#)$CDS: vhdlin version 6.1.8-64b 06/22/2022 16:17 (sjfhw317) $
-- on Mon Dec  2 15:24:48 2024


architecture Structural of nand_2x1 is

begin

    output <= A nand B;

end Structural;
